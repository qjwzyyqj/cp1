module mem_rw_controller;
endmodule
